module ALU_str_1210733 #(parameter n=3)(A , B , Sel , Out)
input signed [n-1:0] A ,B ;
input signed [2:0] Sel ;
output signed reg [n+1:0] ;







endmodule 