module ADD_SUB_1210733#(parameter n=4)(a,b,sel,ans);
input signed [n-1:0]a,b  ; // input size is n
input sel ; // 0 or 1
output reg signed [n:0] ans ; // output size is n+1
always@(a,b,sel)
begin 
	// if the selection is 0 , the block will work as subtracter 
	// and if the selection is 1 , the block will work as adder	
	case(sel)
		1'b0 : ans = a-b ;
		1'b1 : ans = a+b ;
	endcase ;
end
endmodule 